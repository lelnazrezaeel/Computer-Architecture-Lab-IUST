----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:30:05 03/02/2022 
-- Design Name: 
-- Module Name:    XOR_GATE - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity XOR_GATE is
	Port ( a : in  STD_LOGIC;
	b : in STD_LOGIC;
	c : out STD_LOGIC);
end XOR_GATE;

architecture Behavioral of XOR_GATE is
signal z : STD_LOGIC;
begin
z <= a xor b;
c <= z;
end Behavioral;

